-----------------------------------------------------------------------------------
--!     @file    aix4_register_interface_test_bench_64_32.vhd
--!     @brief   AXI4_REGISTER_INTERFACE TEST BENCH(AXI4_DATA_WIDTH=64,REGS_DATA_WIDTH=32)
--!     @version 1.9.0
--!     @date    2023/12/21
--!     @author  Ichiro Kawazome <ichiro_k@ca2.so-net.ne.jp>
-----------------------------------------------------------------------------------
--
--      Copyright (C) 2012-2023 Ichiro Kawazome
--      All rights reserved.
--
--      Redistribution and use in source and binary forms, with or without
--      modification, are permitted provided that the following conditions
--      are met:
--
--        1. Redistributions of source code must retain the above copyright
--           notice, this list of conditions and the following disclaimer.
--
--        2. Redistributions in binary form must reproduce the above copyright
--           notice, this list of conditions and the following disclaimer in
--           the documentation and/or other materials provided with the
--           distribution.
--
--      THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
--      "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
--      LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
--      A PARTICULAR PURPOSE ARE DISCLAIMED.  IN NO EVENT SHALL THE COPYRIGHT
--      OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
--      SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
--      LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
--      DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
--      THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT 
--      (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
--      OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--
-----------------------------------------------------------------------------------
library ieee;
use     ieee.std_logic_1164.all;
entity  AXI4_REGISTER_INTERFACE_TEST_BENCH_64_32 is
    generic (
        NAME            : STRING  := string'("AXI4_REGS_IF_64_32");
        SCENARIO_FILE   : STRING  := string'("axi4_register_interface_test_bench_64_32.snr");
        PRINT_AXI4_READ : boolean := TRUE;
        PRINT_AXI4_WRITE: boolean := TRUE;
        FINISH_ABORT    : boolean := FALSE
    );
end     AXI4_REGISTER_INTERFACE_TEST_BENCH_64_32;
architecture MODEL of AXI4_REGISTER_INTERFACE_TEST_BENCH_64_32 is
begin
    TB: entity work.AXI4_REGISTER_INTERFACE_TEST_BENCH generic map(
            NAME            => NAME,
            SCENARIO_FILE   => SCENARIO_FILE,
            AXI4_DATA_WIDTH => 64,
            REGS_DATA_WIDTH => 32,
            PRINT_AXI4_READ => PRINT_AXI4_READ,
            PRINT_AXI4_WRITE=> PRINT_AXI4_WRITE,
            FINISH_ABORT    => FINISH_ABORT
    );
end MODEL;
